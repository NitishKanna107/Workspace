module comparator(
    
);

endmodule