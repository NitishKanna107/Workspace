module sync_counter(
    input clk, rst,
    output wire[3:0] 
);

endmodule